`ifndef REQ_NUM
`define REQ_NUM 4
`endif

`ifndef EVENT
`define EVENT
event ev;
`endif